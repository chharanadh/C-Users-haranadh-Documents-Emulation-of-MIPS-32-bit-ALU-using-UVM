`define TEST_CASES 1000
`define UVM_TEST   test_throw_random
`define OPERATION Add