`ifndef DEFS_DONE

`define DEFS_DONE
package top_hvl_pkg;
`timescale 1ns/1ps
`include "/pkgs/mentor/questa/10.3/questasim/verilog_src/uvm-1.1d/src/uvm_macros.svh"
///packages required/////// 
import alu_structure_pkg::*;
import uvm_pkg::*;



`include "uvm_macros.svh"
`include "Test_ALU_Constants.sv"


///////////////////////////////
///Including all UVM Files////



//testcases stimulators

`include "test_throw.svh"
`include "test_throw_random.svh"
`include "test_throw_settled.svh"
`include "test_throw_fixed.svh"

//scoreboard
`include "scoreboard.svh"

`include "driver.svh"

//Monitors
`include "monitor1.svh"
`include "monitor2.svh"

//environment classes

`include "environment.svh"
//uvm_test classes
`include "test_throw_fixed_uv.svh"
`include "test_throw_random_uv.svh"
`include "test_throw_settled_uv.svh"
endpackage

import   top_hvl_pkg::*;
`endif